$display ("Verifworks Pvt Ltd");:
